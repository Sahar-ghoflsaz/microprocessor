--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package MyPackage is
constant n: integer :=8;
--constant add : integer:=1;

end MyPackage;

package body MyPackage is
 
end MyPackage;
